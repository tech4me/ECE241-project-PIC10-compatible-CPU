`ifndef DEFINITION_VH
`define DEFINITION_VH

// The constants for status_register
`define STATUS_C 0
`define STATUS_DC 1
`define STATUS_Z 2

`endif