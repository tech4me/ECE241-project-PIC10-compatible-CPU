// This is part of the ECE241 final project
// Date created: November 21 2016
// This file contains functionalitys that helps to monitor all the registers in the cpu

module cpu_watch();

endmodule